`include "config.svh"
`include "game_config.svh"

module lab_top
# (
    parameter  clk_mhz       = 50,
               pixel_mhz     = 25,


               w_key         = 4,
               w_sw          = 8,
               w_led         = 8,
               w_digit       = 8,
               w_gpio        = 100,

               screen_width  = 640,
               screen_height = 480,

               w_red         = 4,
               w_green       = 4,
               w_blue        = 4,

               w_x           = $clog2 ( screen_width  ),
               w_y           = $clog2 ( screen_height ),

               strobe_to_update_xy_counter_width
                   = $clog2 (clk_mhz * 1000 * 1000) - 6
)
(
    input                        clk,
    input                        slow_clk,
    input                        rst,

    // Keys, switches, LEDs

    input        [w_key   - 1:0] key,
    input        [w_sw    - 1:0] sw,
    output logic [w_led   - 1:0] led,

    // A dynamic seven-segment display

    output logic [          7:0] abcdefgh,
    output logic [w_digit - 1:0] digit,

    // Graphics

    input                        display_on,

    input        [w_x     - 1:0] x,
    input        [w_y     - 1:0] y,

    output logic [w_red   - 1:0] red,
    output logic [w_green - 1:0] green,
    output logic [w_blue  - 1:0] blue,

    // Microphone, sound output and UART

    input        [         23:0] mic,
    output       [         15:0] sound,

    input                        uart_rx,
    output                       uart_tx,

    // General-purpose Input/Output

    inout        [w_gpio  - 1:0] gpio
);

    //------------------------------------------------------------------------

       assign led        = '0;
    //    assign abcdefgh   = '0;
    //    assign digit      = '0;
    // assign red        = '0;
    // assign green      = '0;
    // assign blue       = '0;
       assign sound      = '0;
       assign uart_tx    = '1;

    //------------------------------------------------------------------------

    wire [`GAME_RGB_WIDTH - 1:0] rgb;
    logic [2:0] score;
    logic [2:0] n_lifes;
    logic [2:0] debug;

    game_top
    # (
        .clk_mhz                           (clk_mhz                          ),
        .pixel_mhz                         (pixel_mhz                        ),
        .screen_width                      (screen_width                     ),
        .screen_height                     (screen_height                    ),
        .strobe_to_update_xy_counter_width (strobe_to_update_xy_counter_width)
    )
    i_game_top
    (
        .clk              (   clk                ),
        .rst              (   rst                ),

        .launch_key       ( | key                ),
        .left_right_keys  ( { key [3], key [0] } ),
        .shoot  ( key [1] ),

        .display_on       (   display_on         ),

        .x                (   x                  ),
        .y                (   y                  ),

        .score            ( score                ),
        .n_lifes          ( n_lifes              ),
        .debug            ( debug                ),

        .rgb              (   rgb                )
    );



    localparam frame_left   = screen_width * 3 / 10;
    localparam frame_right  = screen_width * 7 / 10;
    localparam frame_top    = 1;
    localparam frame_bottom = screen_height - 1;

    wire on_frame = ((x == frame_left || x == frame_right - 1)  &&
                     (y >= frame_top  && y < frame_bottom) ||
                     (y == frame_top  || y == frame_bottom - 1) &&
                     (x >= frame_left && x < frame_right)
    );

    always_comb begin
        red   = '0;
        green = '0;
        blue  = '0;

        if (on_frame) begin
            red   = { w_red   { 1'b1 } };
            green = { w_green { 1'b1 } };
            blue  = { w_blue  { 1'b1 } };
        end

        if (rgb != 3'b000) begin
            red   = { w_red   { rgb[2] } };
            green = { w_green { rgb[1] } };
            blue  = { w_blue  { rgb[0] } };
        end
    end

    typedef enum bit [7:0]
    {
        ZERO  = 8'b1111_1100,
        ONE   = 8'b0110_0000,
        TWO   = 8'b1101_1010,
        THREE = 8'b1111_0010,
        FOUR  = 8'b0110_0110,
        SPACE = 8'b0000_0000,
        S     = 8'b1011_0110,
        L     = 8'b0001_1100
    }
    seven_seg_encoding_e;

    // logic [3:0] d_digit;
    // always_ff @(posedge clk) begin
    //     if (rst)
    //         d_digit <= 4'b0001;
    //     else
    //         d_digit <= {d_digit[2:0], d_digit[3]};
    // end

    // assign digit = {4'b0000, d_digit};

    // always_comb begin
    //     case (digit)
    //         8'b00000001: abcdefgh = (debug == 0) ? ZERO : (debug == 1) ? ONE : (debug == 2) ? TWO : (debug == 3) ? THREE : (debug == 4) ? FOUR : SPACE;
    //         8'b00000010: abcdefgh = S;
    //         8'b00000100: abcdefgh = (score == 0) ? ZERO : (score == 1) ? ONE : (score == 2) ? TWO : (score == 3) ? THREE : (score == 4) ? FOUR : SPACE;
    //         8'b00001000: abcdefgh = L;
    //         default: abcdefgh = SPACE;
    //     endcase
    // end

// logic [3:0] d_digit;       // To store the digit selection
// logic [15:0] counter;       // Counter to control the pause duration
// parameter MAX_COUNT = 16'd5000;  // Set this value to the desired pause duration
//     always_ff @(posedge clk) begin
//     if (rst) begin
//         d_digit <= 4'b0001;    // Reset d_digit
//         counter <= 0;          // Reset counter
//     end else if (counter == MAX_COUNT) begin
//         counter <= 0;
//         d_digit <= {d_digit[2:0], d_digit[3]}; // Rotate d_digit
//     end else begin
//         counter <= counter + 1; // Increment counter to control pause duration
//     end
//     end

//     assign digit = {4'b0000, d_digit}; // Output digit control (may need adjustment based on your requirements)

//     always_comb begin
//     case (digit)
//         8'b00000001: abcdefgh = (debug == 0) ? ZERO : (debug == 1) ? ONE : (debug == 2) ? TWO : (debug == 3) ? THREE : (debug == 4) ? FOUR : SPACE;
//         8'b00000010: abcdefgh = S;
//         8'b00000100: abcdefgh = (score == 0) ? ZERO : (score == 1) ? ONE : (score == 2) ? TWO : (score == 3) ? THREE : (score == 4) ? FOUR : SPACE;
//         8'b00001000: abcdefgh = L;
//         default: abcdefgh = SPACE;
//     endcase
//     end


/// WORKING ONE
    // logic mux_digit_sel;
    // always_ff @(posedge clk) begin
    //     if (rst)
    //         mux_digit_sel <= 0;
    //     else
    //         mux_digit_sel <= ~mux_digit_sel;
    // end

    // always_comb begin
    // if (mux_digit_sel == 0) begin
    //     abcdefgh = (score == 0) ? ZERO : (score == 1) ? ONE : (score == 2) ? TWO : (score == 3) ? THREE : (score == 4) ? FOUR : SPACE;
    //     digit = 4'b0100;  // активируем младший разряд (предположим 0-й)
    // end else begin
    //     abcdefgh = (debug == 0) ? ZERO : (debug == 1) ? ONE : (debug == 2) ? TWO : (debug == 3) ? THREE : (debug == 4) ? FOUR : SPACE;
    //     digit = 4'b0001;  // активируем старший разряд (1-й)
    // end
    // end

// / THE BEST ONE
    logic [15:0] counter;    // Counter to control the pause duration
    logic mux_digit_sel;

    parameter MAX_COUNT = 16'd5000; // Set this to a value that gives you the desired pause duration

    always_ff @(posedge clk) begin
        if (rst) begin
            mux_digit_sel <= 0;
            counter <= 0;
        end else if (counter == MAX_COUNT) begin
            // Reset counter and toggle mux_digit_sel
            counter <= 0;
            mux_digit_sel <= ~mux_digit_sel;
        end else begin
            counter <= counter + 1;
        end
    end

    always_comb begin
        if (mux_digit_sel == 0) begin
            abcdefgh = (score == 0) ? ZERO : (score == 1) ? ONE : (score == 2) ? TWO : (score == 3) ? THREE : (score == 4) ? FOUR : SPACE;
            digit = 4'b0100;  // Activate lower digit (0th)
        end else begin
            abcdefgh = (debug == 0) ? ZERO : (debug == 1) ? ONE : (debug == 2) ? TWO : (debug == 3) ? THREE : (debug == 4) ? FOUR : SPACE;
            digit = 4'b0001;  // Activate upper digit (1st)
        end
    end


    // assign red   = { w_red   { rgb [2] } };
    // assign green = { w_green { rgb [1] } };
    // assign blue  = { w_blue  { rgb [0] } };

endmodule
