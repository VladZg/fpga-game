`include "config.svh"
`include "game_config.svh"

module lab_top
# (
    parameter  clk_mhz       = 50,
               pixel_mhz     = 25,


               w_key         = 4,
               w_sw          = 8,
               w_led         = 8,
               w_digit       = 8,
               w_gpio        = 100,

               screen_width  = 640,
               screen_height = 480,

               w_red         = 4,
               w_green       = 4,
               w_blue        = 4,

               w_x           = $clog2 ( screen_width  ),
               w_y           = $clog2 ( screen_height ),

               strobe_to_update_xy_counter_width
                   = $clog2 (clk_mhz * 1000 * 1000) - 6
)
(
    input                        clk,
    input                        slow_clk,
    input                        rst,

    // Keys, switches, LEDs

    input        [w_key   - 1:0] key,
    input        [w_sw    - 1:0] sw,
    output logic [w_led   - 1:0] led,

    // A dynamic seven-segment display

    output logic [          7:0] abcdefgh,
    output logic [w_digit - 1:0] digit,

    // Graphics

    input                        display_on,

    input        [w_x     - 1:0] x,
    input        [w_y     - 1:0] y,

    output logic [w_red   - 1:0] red,
    output logic [w_green - 1:0] green,
    output logic [w_blue  - 1:0] blue,

    // Microphone, sound output and UART

    input        [         23:0] mic,
    output       [         15:0] sound,

    input                        uart_rx,
    output                       uart_tx,

    // General-purpose Input/Output

    inout        [w_gpio  - 1:0] gpio
);

    //------------------------------------------------------------------------

       assign led        = '0;
       assign abcdefgh   = '0;
       assign digit      = '0;
    // assign red        = '0;
    // assign green      = '0;
    // assign blue       = '0;
       assign sound      = '0;
       assign uart_tx    = '1;

    //------------------------------------------------------------------------

    wire [`GAME_RGB_WIDTH - 1:0] rgb;

    game_top
    # (
        .clk_mhz                           (clk_mhz                          ),
        .pixel_mhz                         (pixel_mhz                        ),
        .screen_width                      (screen_width                     ),
        .screen_height                     (screen_height                    ),
        .strobe_to_update_xy_counter_width (strobe_to_update_xy_counter_width)
    )
    i_game_top
    (
        .clk              (   clk                ),
        .rst              (   rst                ),

        .launch_key       ( | key                ),
        .left_right_keys  ( { key [3], key [0] } ),
        .shoot  ( key [1] ),

        .display_on       (   display_on         ),

        .x                (   x                  ),
        .y                (   y                  ),

        .rgb              (   rgb                )
    );


    logic [63:0] sprite [0:15] = '{
        64'h0000000000000000,
        64'h0000000000ff0ff0,
        64'h000000000fccfc90,
        64'h000000000fccccbf,
        64'h00fff000fffcccf0,
        64'h0fcccf0fcccfcf00,
        64'hfcccccfccbbcf000,
        64'hfcccccccccbcf000,
        64'hfcccccccccccf000,
        64'h0fcccccccccf0000,
        64'h00fcccccccf00000,
        64'h000fcccccf000000,
        64'h0000fcccf0000000,
        64'h00000fcf00000000,
        64'h000000f000000000,
        64'h0000000000000000
    };

    // --- Спрайт 16×16 в левом верхнем углу (используем младшие 16 бит каждой строки) ---
    logic [63:0] sprite [0:15] = '{
        64'h0000000000000000,
        64'h0000000000ff0ff0,
        64'h000000000fccfc90,
        64'h000000000fccccbf,
        64'h00fff000fffcccf0,
        64'h0fcccf0fcccfcf00,
        64'hfcccccfccbbcf000,
        64'hfcccccccccbcf000,
        64'hfcccccccccccf000,
        64'h0fcccccccccf0000,
        64'h00fcccccccf00000,
        64'h000fcccccf000000,
        64'h0000fcccf0000000,
        64'h00000fcf00000000,
        64'h000000f000000000,
        64'h0000000000000000
    };

    wire in_sprite_bounds  = (x < 16) && (y < 16);
    wire sprite_pixel_on   = in_sprite_bounds && sprite[y][63 - x];

    localparam frame_left   = screen_width  / 4;
    localparam frame_right  = screen_width  * 3 / 4;
    localparam frame_top    = screen_height / 4;
    localparam frame_bottom = screen_height * 3 / 4;

    wire on_frame = (
           (x == frame_left  || x == frame_right - 1) && (y >= frame_top && y < frame_bottom)
        || (y == frame_top   || y == frame_bottom - 1) && (x >= frame_left && x < frame_right)
    );

    always_comb begin
        red   = '0;
        green = '0;
        blue  = '0;

        if (on_frame) begin
            red   = { w_red   { 1'b1 } };
            green = { w_green { 1'b1 } };
            blue  = { w_blue  { 1'b1 } };
        end

        if (sprite_pixel_on) begin
            red   = { w_red   { 1'b1 } };
            green = { w_green { 1'b1 } };
            blue  = { w_blue  { 1'b1 } };
        end

        if (rgb != 3'b000) begin
            red   = { w_red   { rgb[2] } };
            green = { w_green { rgb[1] } };
            blue  = { w_blue  { rgb[0] } };
        end
    end



    // assign red   = { w_red   { rgb [2] } };
    // assign green = { w_green { rgb [1] } };
    // assign blue  = { w_blue  { rgb [0] } };

endmodule
